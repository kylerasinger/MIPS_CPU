
-- set up vcom source
source /CMC/ENVIRONMENT/modelsim.env


-- set up xilinx source
source /CMC/tools/xilinx/Vivado_2018.2/Vivado/2018.2/settings64_CMC_central_license.csh
