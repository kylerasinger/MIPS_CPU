library IEEE;
use IEEE.std_logic_1164.all;
--use IEEE.numeric_std.all;
use IEEE.std_logic_signed.all;

entity next_address is
	port(
		rt, rs : in std_logic_vector(31 downto 0); 			-- two register inputs (defined in opcode)
		pc : in std_logic_vector(31 downto 0);				-- PC register
		target_address : in std_logic_vector(25 downto 0);	-- address to jump to (can be bottom 16)
		branch_type : in std_logic_vector(1 downto 0);		-- type of branch (generated by control unit)
			-- 00 is non branch instructions
			-- 01 is beq instr.
			-- 10 is bne instr.
			-- 11 is bltz
		pc_sel : in std_logic_vector(1 downto 0);			-- type of jump(generated by control unit)
			-- 00 is non jump instructions
			-- 01 is jump instructions
			-- 10 is jump register instructions
			-- 11 unused

		next_pc : out std_logic_vector(31 downto 0)			-- the next PC position in execution
	);	
end next_address ;

architecture my_next_address of next_address is

	signal temp_pc : std_logic_vector(31 downto 0);

begin

	process(rt, rs, pc, target_address, branch_type, pc_sel, temp_pc)
	
	begin
		
		-- Branch type logic
		case branch_type is
			when "00" =>
				-- no branch
				temp_pc <= std_logic_vector((pc) + X"00000001");
			when "01" =>
				-- beq instruction (branch if equal)
				if (rs /= rt) then
					temp_pc <= std_logic_vector((pc) + X"00000001");
				else
					-- sign extension for the other 16 bits
					temp_pc <= pc + X"00000001" + ((31 downto 16 => target_address(15)) & target_address(15 downto 0));					
				end if;
			when "10" =>
				-- bne (branch not equal)
				if (rs /= rt) then
					temp_pc <= pc + 1 + ((31 downto 16 => target_address(15)) & target_address(15 downto 0));
				else
					temp_pc <= std_logic_vector((pc) + X"00000001");

				end if;
			when "11" =>
				-- bltz (branch less than zero AKA, branch if rs is negative)
				if (rs(31) = '1') then
					temp_pc <= pc + 1 + ((31 downto 16 => target_address(15)) & target_address(15 downto 0));
				else
					temp_pc <= std_logic_vector((pc) + X"00000001");

				end if;	
			when others =>
				temp_pc <= std_logic_vector((pc) + X"00000001");
		end case;

		-- PC selection logic
		case pc_sel is
		    when "00" =>
		        next_pc <= temp_pc;  -- select compute next pc, must be =00 for branch type
		    when "01" =>
		        next_pc <= "000000" & target_address(25 downto 0);  -- Jump to target address
		    when "10" =>
		        next_pc <= rs;  -- next PC is the register source
		    when others =>
		        next_pc <= pc;  -- not used
		end case;

	end process;
end my_next_address;
































