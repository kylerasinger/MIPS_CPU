library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_signed.all;

entity cpu is
	port(
		-- I changed the names of the signals, must change in the XDC and .do
		reset		: in std_logic;
		clk		: in std_logic;

		rs_out, rt_out	: out std_logic_vector(3 downto 0) := (others => '0');
		pc_out		: out std_logic_vector(3 downto 0) := (others => '0');
		overflow, zero	: out std_logic
	);
end cpu;

architecture my_cpu of cpu is
	
	-----= Start of Component Declaration =------
	
	-- lab 1
	component alu
		port(
			-- IN
			x, y 		: in std_logic_vector(31 downto 0);
			add_sub 	: in std_logic ; 
					-- 0 = add, 1 = sub
			logic_func 	: in std_logic_vector(1 downto 0) ;
					-- 00 AND, 01 OR, 10 XOR, 11 NOR
			func 		: in std_logic_vector(1 downto 0) ; 
					-- 00 = lui, 01 = setless, 10 = arith, 11 = logic
			-- OUT
			output 		: out std_logic_vector(31 downto 0);
			overflow 	: out std_logic;
			zero 		: out std_logic 
		); 
	end component;

	-- lab 2
	component regfile
		port( 
			-- IN
			din 		: in std_logic_vector(31 downto 0);				
					--data to be written
			reg_reset 		: in std_logic; 	
					--sets all to 0 when == 1
			clk 		: in std_logic;
			write 		: in std_logic;
					--writes to write_address (sync)
			read_a 		: in std_logic_vector(4 downto 0);			
					--address for out_a reg (async)
			read_b 		: in std_logic_vector(4 downto 0);			
					--address for out_b reg (async)
			write_address 	: in std_logic_vector(4 downto 0);	
					--address for din to be written to (sync)

			-- OUT
			out_a : out std_logic_vector(31 downto 0);
			out_b : out std_logic_vector(31 downto 0)
		);
	end component;

	-- lab 3
	component next_address
		port(
			-- IN
			rt, rs 		: in std_logic_vector(31 downto 0);
					-- two register inputs (defined in opcode)
			pc 		: in std_logic_vector(31 downto 0);
					-- PC register
			target_address 	: in std_logic_vector(25 downto 0);
					-- address to jump to (can be bottom 16)
			branch_type 	: in std_logic_vector(1 downto 0);
					-- type of branch (generated by control unit)
						-- 00 is non branch instructions
						-- 01 is beq instr.
						-- 10 is bne instr.
						-- 11 is bltz
			pc_sel 		: in std_logic_vector(1 downto 0);
					-- type of jump(generated by control unit)
						-- 00 is non jump instructions
						-- 01 is jump instructions
						-- 10 is jump register instructions
						-- 11 unused
			-- OUT
			next_pc 	: out std_logic_vector(31 downto 0)			
					-- the next PC position in execution
		);	
	end component;

	--lab 4 onwards
	component pc_register
		port(
			pc_in 		: in std_logic_vector(31 downto 0);
			pc_reset 	: in std_logic;
			clk		: in std_logic;
			
			pc_out 		: out std_logic_vector(31 downto 0)
		);
	end component;

	component ic_cache
		port(
			address		: in std_logic_vector(4 downto 0);
			
			instruction	: out std_logic_vector(31 downto 0)
		);
	end component;

	component data_cache
		port(
			data_in		: in std_logic_vector(31 downto 0);
		    	dc_reset     	: in std_logic;
		    	clk       	: in std_logic;
		    	address  	: in std_logic_vector(4 downto 0);
		    	data_write	: in std_logic;
	 
		    	data_out     	: out std_logic_vector(31 downto 0)
		);
	end component;

	component sign_extender
		port(
			input		: in std_logic_vector(15 downto 0);
			func    	: in std_logic_vector(1 downto 0);

			output 		: out std_logic_vector(31 downto 0)
		);
	end component;
	
	-----=  End of Component Declaration  =------

	-- Component Configuration
	for a_alu 		: alu use entity WORK.alu(my_alu);
	for a_regfile		: regfile use entity WORK.regfile(my_regfile);
	for a_next_address	: next_address use entity WORK.next_address(my_next_address);
	for a_pc_register	: pc_register use entity WORK.pc_register(my_pc_register);
	for a_ic_cache		: ic_cache use entity WORK.ic_cache(my_ic_cache);
	for a_data_cache	: data_cache use entity WORK.data_cache(my_data_cache);
	for a_sign_extender	: sign_extender use entity WORK.sign_extender(my_sign_extender);

	-----= Start of Databus Signals =-----

	-- Component Outputs
		-- ALU
		signal alu_out 			: std_logic_vector(31 downto 0) := X"00000000";
		-- REGFILE
		signal reg_out_a, reg_out_b	: std_logic_vector(31 downto 0) := X"00000000";
		-- NEXT ADDRESS
		signal next_pc_out 		: std_logic_vector(31 downto 0) := X"00000000";
		-- PC REGISTER
		signal pc_reg_out	 	: std_logic_vector(31 downto 0) := X"00000000";
		-- I CACHE
		signal i_cache_out 		: std_logic_vector(31 downto 0) := X"00000000";
		-- D CACHE
		signal data_cache_out 		: std_logic_vector(31 downto 0) := X"00000000";
		-- SIGN EXTENDER
		signal sign_ext_out 		: std_logic_vector(31 downto 0) := X"00000000";
	-- Split Signals
	-- Control Unit Signals
		signal c_reg_write 		: std_logic := '0';
		signal c_add_sub 		: std_logic := '0';
		signal c_logic_func, c_func	: std_logic_vector(1 downto 0) := "00";
		signal c_branch_type, c_pc_sel	: std_logic_vector(1 downto 0) := "00";
		signal c_data_write		: std_logic := '0';
		signal cc_opcode, cc_func	: std_logic_vector(5 downto 0) := "000000";
		signal cc_control_signal	: std_logic_vector(11 downto 0) := "000000000000";
	-- Mux Signals
		signal reg_dst, alu_src, reg_in_src : std_logic := '0';
		signal mux1_out 		: std_logic_vector(4 downto 0) := "00000";
		signal mux2_out 		: std_logic_vector(31 downto 0) := X"00000000";
		signal mux3_out 		: std_logic_vector(31 downto 0) := X"00000000";

	-----=  End of Databus Signals  =-----

	begin

	-----= Start of Control Unit =-----

	process(clk, i_cache_out, reset, cc_opcode, cc_func, cc_control_signal)
	begin
		cc_opcode <= i_cache_out(31 downto 26);
		cc_func <= i_cache_out(5 downto 0);
		cc_control_signal <= cc_opcode & cc_func;
		
		case cc_opcode is
			-- lui
			when "001111" =>
				c_reg_write <= 		'1';
				reg_dst <= 		'0';
				reg_in_src <= 		'1';
				alu_src <= 		'1';
				c_add_sub <= 		'0';
				c_data_write <= 	'0';
				c_logic_func <= 	"00";
				c_func <= 		"00";
				c_branch_type <=	"00";
				c_pc_sel <=		"00";
			-- ALU
			when "000000" =>
				-- add
				if cc_func = "100000" then
					c_reg_write <= 		'1';
					reg_dst <= 		'1';
					reg_in_src <= 		'1';
					alu_src <= 		'0';
					c_add_sub <= 		'0';
					c_data_write <= 	'0';
					c_logic_func <= 	"00";
					c_func <= 		"10";
					c_branch_type <=	"00";
					c_pc_sel <=		"00";
				-- sub
				elsif cc_func = "100010" then 
					c_reg_write <= 		'1';
					reg_dst <= 		'1';
					reg_in_src <= 		'1';
					alu_src <= 		'0';
					c_add_sub <= 		'1';
					c_data_write <= 	'0';
					c_logic_func <= 	"00";
					c_func <= 		"10";
					c_branch_type <=	"00";
					c_pc_sel <=		"00";
				-- slt
				elsif cc_func = "101010" then
					c_reg_write <= 		'1';
					reg_dst <= 		'1';
					reg_in_src <= 		'1';
					alu_src <= 		'0';
					c_add_sub <= 		'1';
					c_data_write <= 	'0';
					c_logic_func <= 	"00";
					c_func <= 		"01";
					c_branch_type <=	"00";
					c_pc_sel <=		"00";
				-- and	
				elsif cc_func = "100100" then
					c_reg_write <= 		'1';
					reg_dst <= 		'1';
					reg_in_src <= 		'1';
					alu_src <= 		'0';
					c_add_sub <= 		'1';
					c_data_write <= 	'0';
					c_logic_func <= 	"00";
					c_func <= 		"11";
					c_branch_type <=	"00";
					c_pc_sel <=		"00";
				-- or
				elsif cc_func = "100101" then
					c_reg_write <= 		'1';
					reg_dst <= 		'1';
					reg_in_src <= 		'1';
					alu_src <= 		'0';
					c_add_sub <= 		'1';
					c_data_write <= 	'0';
					c_logic_func <= 	"01";
					c_func <= 		"11";
					c_branch_type <=	"00";
					c_pc_sel <=		"00";
				-- xor
				elsif cc_func = "100110" then
					c_reg_write <= 		'1';
					reg_dst <= 		'1';
					reg_in_src <= 		'1';
					alu_src <= 		'0';
					c_add_sub <= 		'1';
					c_data_write <= 	'0';
					c_logic_func <= 	"10";
					c_func <= 		"11";
					c_branch_type <=	"00";
					c_pc_sel <=		"00";
				-- nor
				elsif cc_func = "100111" then
					c_reg_write <= 		'1';
					reg_dst <= 		'1';
					reg_in_src <= 		'1';
					alu_src <= 		'0';
					c_add_sub <= 		'1';
					c_data_write <= 	'0';
					c_logic_func <= 	"11";
					c_func <= 		"11";
					c_branch_type <=	"00";
					c_pc_sel <=		"00";
				-- jr
				elsif cc_func = "001000" then
					c_reg_write <= 		'0';
					reg_dst <= 		'0';
					reg_in_src <= 		'0';
					alu_src <= 		'0';
					c_add_sub <= 		'0';
					c_data_write <= 	'0';
					c_logic_func <= 	"00";
					c_func <= 		"00";
					c_branch_type <=	"00";
					c_pc_sel <=		"10";			
				end if;

			-- addi
			when "001000" =>
				c_reg_write <= 		'1';
				reg_dst <= 		'0';
				reg_in_src <= 		'1';
				alu_src <= 		'1';
				c_add_sub <= 		'0';
				c_data_write <= 	'0';
				c_logic_func <= 	"00";
				c_func <= 		"10";
				c_branch_type <=	"00";
				c_pc_sel <=		"00";
			-- slti
			when "001010" =>
				c_reg_write <= 		'1';
				reg_dst <= 		'0';
				reg_in_src <= 		'1';
				alu_src <= 		'1';
				c_add_sub <= 		'1';
				c_data_write <= 	'0';
				c_logic_func <= 	"00";
				c_func <= 		"01";
				c_branch_type <=	"00";
				c_pc_sel <=		"00";
			-- andi
			when "001100" =>
				c_reg_write <= 		'1';
				reg_dst <= 		'0';
				reg_in_src <= 		'1';
				alu_src <= 		'1';
				c_add_sub <= 		'1';
				c_data_write <= 	'0';
				c_logic_func <= 	"00";
				c_func <= 		"11";
				c_branch_type <=	"00";
				c_pc_sel <=		"00";
			-- ori
			when "001101" =>
				c_reg_write <= 		'1';
				reg_dst <= 		'0';
				reg_in_src <= 		'1';
				alu_src <= 		'1';
				c_add_sub <= 		'1';
				c_data_write <= 	'0';
				c_logic_func <= 	"01";
				c_func <= 		"11";
				c_branch_type <=	"00";
				c_pc_sel <=		"00";
			-- xori
			when "001110" =>
				c_reg_write <= 		'1';
				reg_dst <= 		'0';
				reg_in_src <= 		'1';
				alu_src <= 		'1';
				c_add_sub <= 		'1';
				c_data_write <= 	'0';
				c_logic_func <= 	"10";
				c_func <= 		"11";
				c_branch_type <=	"00";
				c_pc_sel <=		"00";
			-- lw
			when "100011" =>
				c_reg_write <= 		'1';
				reg_dst <= 		'0';
				reg_in_src <= 		'0';
				alu_src <= 		'1';
				c_add_sub <= 		'0';
				c_data_write <= 	'0';
				c_logic_func <= 	"10";
				c_func <= 		"10";
				c_branch_type <=	"00";
				c_pc_sel <=		"00";
			-- sw
			when "101011" =>
				c_reg_write <= 		'0';
				reg_dst <= 		'0';
				reg_in_src <= 		'0';
				alu_src <= 		'1';
				c_add_sub <= 		'0';
				c_data_write <= 	'1';
				c_logic_func <= 	"10";
				c_func <= 		"10";
				c_branch_type <=	"00";
				c_pc_sel <=		"00";
			-- j
			when "000010" =>
				c_reg_write <= 		'0';
				reg_dst <= 		'0';
				reg_in_src <= 		'0';
				alu_src <= 		'0';
				c_add_sub <= 		'0';
				c_data_write <= 	'0';
				c_logic_func <= 	"00";
				c_func <= 		"00";
				c_branch_type <=	"00";
				c_pc_sel <=		"01";
			-- bltz
			when "000001" =>
				c_reg_write <= 		'0';
				reg_dst <= 		'0';
				reg_in_src <= 		'0';
				alu_src <= 		'0';
				c_add_sub <= 		'0';
				c_data_write <= 	'0';
				c_logic_func <= 	"00";
				c_func <= 		"00";
				c_branch_type <=	"11";
				c_pc_sel <=		"00";
			-- beq
			when "000100" =>
				c_reg_write <= 		'0';
				reg_dst <= 		'0';
				reg_in_src <= 		'0';
				alu_src <= 		'0';
				c_add_sub <= 		'0';
				c_data_write <= 	'0';
				c_logic_func <= 	"00";
				c_func <= 		"00";
				c_branch_type <=	"01";
				c_pc_sel <=		"00";
			-- bne
			when "000101" =>
				c_reg_write <= 		'0';
				reg_dst <= 		'0';
				reg_in_src <= 		'0';
				alu_src <= 		'0';
				c_add_sub <= 		'0';
				c_data_write <= 	'0';
				c_logic_func <= 	"00";
				c_func <= 		"00";
				c_branch_type <=	"10";
				c_pc_sel <=		"00";
			when others =>
				c_reg_write <= '0';
			
		
		end case;	
			
	end process;
	-----=  End of Control Unit  =-----

	-----= Start of Component Instantiation =------

	a_alu: alu port map(
		--in		
			x => reg_out_a,
			y => mux2_out,
			add_sub => c_add_sub,
			logic_func => c_logic_func,
			func => c_func,
		--out
			output => alu_out,
			overflow => overflow,
			zero => zero
	);

	a_regfile: regfile port map(
		-- in
			din => mux3_out,
			reg_reset => reset,
			clk => clk,		
			write => c_reg_write,
			read_a => i_cache_out(25 downto 21),
			read_b => i_cache_out(20 downto 16),
			write_address => mux1_out,
		-- out
			out_a => reg_out_a,
			out_b => reg_out_b
	);
	
	a_next_address: next_address port map(
		-- in
			rt => reg_out_a, 
			rs => reg_out_b,
			pc => pc_reg_out,
			target_address => i_cache_out(25 downto 0),
			branch_type => c_branch_type,
			pc_sel => c_pc_sel,
		-- out
			next_pc => next_pc_out
	);

	a_pc_register: pc_register port map(
		-- in			
			pc_in => next_pc_out,
			pc_reset => reset,
			clk => clk,
		-- out
			pc_out => pc_reg_out
	);

	a_ic_cache: ic_cache port map(
		-- in
			address => pc_reg_out(4 downto 0),
		-- out
			instruction => i_cache_out
	);

	a_data_cache: data_cache port map(
		-- in
			data_in => reg_out_b,
		    	dc_reset => reset,
		    	clk => clk,
		    	address => alu_out(4 downto 0),
		    	data_write => c_data_write,
		-- out
		    	data_out => data_cache_out
	);

	a_sign_extender: sign_extender port map(
		-- in
			input => i_cache_out(15 downto 0),
			func => c_func,
		-- out
			output => sign_ext_out
	);
	
	-----=  End of Component Instantiation  =------

	-----= Start of Multiplexers =-----

		-- Mux 1
		mux1_out <= 
			i_cache_out(20 downto 16) when (reg_dst = '0') else
			i_cache_out(15 downto 11) when (reg_dst = '1');
				
		-- Mux 2
		mux2_out <=
			reg_out_b(31 downto 0) when (alu_src = '0') else
			sign_ext_out(31 downto 0) when (alu_src = '1');

		-- Mux 3
		mux3_out <=
			data_cache_out(31 downto 0) when (reg_in_src = '0') else
			alu_out(31 downto 0) when (reg_in_src = '1');

	-----=  End of Multiplexers  =-----

	rs_out <= reg_out_a(3 downto 0);
	rt_out <= reg_out_b(3 downto 0);
	pc_out <= pc_reg_out(3 downto 0);

end my_cpu;
	

